
module onchipAlarm (
	clk_clk,
	reset_reset_n,
	led_export);	

	input		clk_clk;
	input		reset_reset_n;
	output		led_export;
endmodule
