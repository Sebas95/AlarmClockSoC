
module onchipAlarm (
	clk_clk,
	led_export,
	reset_reset_n);	

	input		clk_clk;
	output		led_export;
	input		reset_reset_n;
endmodule
