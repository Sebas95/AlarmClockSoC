// onchipAlarm.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module onchipAlarm (
		input  wire       clk_clk,             //          clk.clk
		output wire [6:0] horas_d_export,      //      horas_d.export
		output wire [6:0] horas_u_export,      //      horas_u.export
		output wire       led_export,          //          led.export
		output wire [6:0] minutos_d_export,    //    minutos_d.export
		output wire [6:0] minutos_u_export,    //    minutos_u.export
		input  wire       modo_export,         //         modo.export
		input  wire [3:0] push_buttons_export, // push_buttons.export
		input  wire       reset_reset_n,       //        reset.reset_n
		output wire [6:0] segundos_d_export,   //   segundos_d.export
		output wire [6:0] segundos_u_export    //   segundos_u.export
	);

	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [15:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [15:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [11:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_led_s1_chipselect;                         // mm_interconnect_0:led_s1_chipselect -> led:chipselect
	wire  [31:0] mm_interconnect_0_led_s1_readdata;                           // led:readdata -> mm_interconnect_0:led_s1_readdata
	wire   [1:0] mm_interconnect_0_led_s1_address;                            // mm_interconnect_0:led_s1_address -> led:address
	wire         mm_interconnect_0_led_s1_write;                              // mm_interconnect_0:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_0_led_s1_writedata;                          // mm_interconnect_0:led_s1_writedata -> led:writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                     // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                       // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                        // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                          // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                      // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire  [31:0] mm_interconnect_0_push_buttons_s1_readdata;                  // push_buttons:readdata -> mm_interconnect_0:push_buttons_s1_readdata
	wire   [1:0] mm_interconnect_0_push_buttons_s1_address;                   // mm_interconnect_0:push_buttons_s1_address -> push_buttons:address
	wire  [31:0] mm_interconnect_0_modo_s1_readdata;                          // modo:readdata -> mm_interconnect_0:modo_s1_readdata
	wire   [1:0] mm_interconnect_0_modo_s1_address;                           // mm_interconnect_0:modo_s1_address -> modo:address
	wire         mm_interconnect_0_horas_d_s1_chipselect;                     // mm_interconnect_0:horas_d_s1_chipselect -> horas_d:chipselect
	wire  [31:0] mm_interconnect_0_horas_d_s1_readdata;                       // horas_d:readdata -> mm_interconnect_0:horas_d_s1_readdata
	wire   [1:0] mm_interconnect_0_horas_d_s1_address;                        // mm_interconnect_0:horas_d_s1_address -> horas_d:address
	wire         mm_interconnect_0_horas_d_s1_write;                          // mm_interconnect_0:horas_d_s1_write -> horas_d:write_n
	wire  [31:0] mm_interconnect_0_horas_d_s1_writedata;                      // mm_interconnect_0:horas_d_s1_writedata -> horas_d:writedata
	wire         mm_interconnect_0_horas_u_s1_chipselect;                     // mm_interconnect_0:horas_u_s1_chipselect -> horas_u:chipselect
	wire  [31:0] mm_interconnect_0_horas_u_s1_readdata;                       // horas_u:readdata -> mm_interconnect_0:horas_u_s1_readdata
	wire   [1:0] mm_interconnect_0_horas_u_s1_address;                        // mm_interconnect_0:horas_u_s1_address -> horas_u:address
	wire         mm_interconnect_0_horas_u_s1_write;                          // mm_interconnect_0:horas_u_s1_write -> horas_u:write_n
	wire  [31:0] mm_interconnect_0_horas_u_s1_writedata;                      // mm_interconnect_0:horas_u_s1_writedata -> horas_u:writedata
	wire         mm_interconnect_0_minutos_d_s1_chipselect;                   // mm_interconnect_0:minutos_d_s1_chipselect -> minutos_d:chipselect
	wire  [31:0] mm_interconnect_0_minutos_d_s1_readdata;                     // minutos_d:readdata -> mm_interconnect_0:minutos_d_s1_readdata
	wire   [1:0] mm_interconnect_0_minutos_d_s1_address;                      // mm_interconnect_0:minutos_d_s1_address -> minutos_d:address
	wire         mm_interconnect_0_minutos_d_s1_write;                        // mm_interconnect_0:minutos_d_s1_write -> minutos_d:write_n
	wire  [31:0] mm_interconnect_0_minutos_d_s1_writedata;                    // mm_interconnect_0:minutos_d_s1_writedata -> minutos_d:writedata
	wire         mm_interconnect_0_minutos_u_s1_chipselect;                   // mm_interconnect_0:minutos_u_s1_chipselect -> minutos_u:chipselect
	wire  [31:0] mm_interconnect_0_minutos_u_s1_readdata;                     // minutos_u:readdata -> mm_interconnect_0:minutos_u_s1_readdata
	wire   [1:0] mm_interconnect_0_minutos_u_s1_address;                      // mm_interconnect_0:minutos_u_s1_address -> minutos_u:address
	wire         mm_interconnect_0_minutos_u_s1_write;                        // mm_interconnect_0:minutos_u_s1_write -> minutos_u:write_n
	wire  [31:0] mm_interconnect_0_minutos_u_s1_writedata;                    // mm_interconnect_0:minutos_u_s1_writedata -> minutos_u:writedata
	wire         mm_interconnect_0_segundos_u_s1_chipselect;                  // mm_interconnect_0:segundos_u_s1_chipselect -> segundos_u:chipselect
	wire  [31:0] mm_interconnect_0_segundos_u_s1_readdata;                    // segundos_u:readdata -> mm_interconnect_0:segundos_u_s1_readdata
	wire   [1:0] mm_interconnect_0_segundos_u_s1_address;                     // mm_interconnect_0:segundos_u_s1_address -> segundos_u:address
	wire         mm_interconnect_0_segundos_u_s1_write;                       // mm_interconnect_0:segundos_u_s1_write -> segundos_u:write_n
	wire  [31:0] mm_interconnect_0_segundos_u_s1_writedata;                   // mm_interconnect_0:segundos_u_s1_writedata -> segundos_u:writedata
	wire         mm_interconnect_0_segundos_d_s1_chipselect;                  // mm_interconnect_0:segundos_d_s1_chipselect -> segundos_d:chipselect
	wire  [31:0] mm_interconnect_0_segundos_d_s1_readdata;                    // segundos_d:readdata -> mm_interconnect_0:segundos_d_s1_readdata
	wire   [1:0] mm_interconnect_0_segundos_d_s1_address;                     // mm_interconnect_0:segundos_d_s1_address -> segundos_d:address
	wire         mm_interconnect_0_segundos_d_s1_write;                       // mm_interconnect_0:segundos_d_s1_write -> segundos_d:write_n
	wire  [31:0] mm_interconnect_0_segundos_d_s1_writedata;                   // mm_interconnect_0:segundos_d_s1_writedata -> segundos_d:writedata
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // timer_0:irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [horas_d:reset_n, horas_u:reset_n, led:reset_n, minutos_d:reset_n, minutos_u:reset_n, mm_interconnect_0:led_reset_reset_bridge_in_reset_reset, modo:reset_n, push_buttons:reset_n, segundos_d:reset_n, segundos_u:reset_n, timer_0:reset_n]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_memory2_0:reset, rst_translator:in_reset]
	wire         rst_controller_001_reset_out_reset_req;                      // rst_controller_001:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                      // nios2_gen2_0:debug_reset_request -> rst_controller_001:reset_in1

	onchipAlarm_horas_d horas_d (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_horas_d_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_horas_d_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_horas_d_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_horas_d_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_horas_d_s1_readdata),   //                    .readdata
		.out_port   (horas_d_export)                           // external_connection.export
	);

	onchipAlarm_horas_d horas_u (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_horas_u_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_horas_u_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_horas_u_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_horas_u_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_horas_u_s1_readdata),   //                    .readdata
		.out_port   (horas_u_export)                           // external_connection.export
	);

	onchipAlarm_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	onchipAlarm_led led (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (led_export)                           // external_connection.export
	);

	onchipAlarm_horas_d minutos_d (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_minutos_d_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_minutos_d_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_minutos_d_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_minutos_d_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_minutos_d_s1_readdata),   //                    .readdata
		.out_port   (minutos_d_export)                           // external_connection.export
	);

	onchipAlarm_horas_d minutos_u (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_minutos_u_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_minutos_u_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_minutos_u_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_minutos_u_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_minutos_u_s1_readdata),   //                    .readdata
		.out_port   (minutos_u_export)                           // external_connection.export
	);

	onchipAlarm_modo modo (
		.clk      (clk_clk),                            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address  (mm_interconnect_0_modo_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_modo_s1_readdata), //                    .readdata
		.in_port  (modo_export)                         // external_connection.export
	);

	onchipAlarm_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	onchipAlarm_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),           //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	onchipAlarm_push_buttons push_buttons (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_push_buttons_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_push_buttons_s1_readdata), //                    .readdata
		.in_port  (push_buttons_export)                         // external_connection.export
	);

	onchipAlarm_horas_d segundos_d (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_segundos_d_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_segundos_d_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_segundos_d_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_segundos_d_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_segundos_d_s1_readdata),   //                    .readdata
		.out_port   (segundos_d_export)                           // external_connection.export
	);

	onchipAlarm_horas_d segundos_u (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_segundos_u_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_segundos_u_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_segundos_u_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_segundos_u_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_segundos_u_s1_readdata),   //                    .readdata
		.out_port   (segundos_u_export)                           // external_connection.export
	);

	onchipAlarm_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	onchipAlarm_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                     //                                clk_0_clk.clk
		.led_reset_reset_bridge_in_reset_reset          (rst_controller_reset_out_reset),                              //          led_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                            //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                        //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                         //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                               //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                           //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                              //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                          //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                        //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                     //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                 //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                        //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                    //                                         .readdata
		.horas_d_s1_address                             (mm_interconnect_0_horas_d_s1_address),                        //                               horas_d_s1.address
		.horas_d_s1_write                               (mm_interconnect_0_horas_d_s1_write),                          //                                         .write
		.horas_d_s1_readdata                            (mm_interconnect_0_horas_d_s1_readdata),                       //                                         .readdata
		.horas_d_s1_writedata                           (mm_interconnect_0_horas_d_s1_writedata),                      //                                         .writedata
		.horas_d_s1_chipselect                          (mm_interconnect_0_horas_d_s1_chipselect),                     //                                         .chipselect
		.horas_u_s1_address                             (mm_interconnect_0_horas_u_s1_address),                        //                               horas_u_s1.address
		.horas_u_s1_write                               (mm_interconnect_0_horas_u_s1_write),                          //                                         .write
		.horas_u_s1_readdata                            (mm_interconnect_0_horas_u_s1_readdata),                       //                                         .readdata
		.horas_u_s1_writedata                           (mm_interconnect_0_horas_u_s1_writedata),                      //                                         .writedata
		.horas_u_s1_chipselect                          (mm_interconnect_0_horas_u_s1_chipselect),                     //                                         .chipselect
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.led_s1_address                                 (mm_interconnect_0_led_s1_address),                            //                                   led_s1.address
		.led_s1_write                                   (mm_interconnect_0_led_s1_write),                              //                                         .write
		.led_s1_readdata                                (mm_interconnect_0_led_s1_readdata),                           //                                         .readdata
		.led_s1_writedata                               (mm_interconnect_0_led_s1_writedata),                          //                                         .writedata
		.led_s1_chipselect                              (mm_interconnect_0_led_s1_chipselect),                         //                                         .chipselect
		.minutos_d_s1_address                           (mm_interconnect_0_minutos_d_s1_address),                      //                             minutos_d_s1.address
		.minutos_d_s1_write                             (mm_interconnect_0_minutos_d_s1_write),                        //                                         .write
		.minutos_d_s1_readdata                          (mm_interconnect_0_minutos_d_s1_readdata),                     //                                         .readdata
		.minutos_d_s1_writedata                         (mm_interconnect_0_minutos_d_s1_writedata),                    //                                         .writedata
		.minutos_d_s1_chipselect                        (mm_interconnect_0_minutos_d_s1_chipselect),                   //                                         .chipselect
		.minutos_u_s1_address                           (mm_interconnect_0_minutos_u_s1_address),                      //                             minutos_u_s1.address
		.minutos_u_s1_write                             (mm_interconnect_0_minutos_u_s1_write),                        //                                         .write
		.minutos_u_s1_readdata                          (mm_interconnect_0_minutos_u_s1_readdata),                     //                                         .readdata
		.minutos_u_s1_writedata                         (mm_interconnect_0_minutos_u_s1_writedata),                    //                                         .writedata
		.minutos_u_s1_chipselect                        (mm_interconnect_0_minutos_u_s1_chipselect),                   //                                         .chipselect
		.modo_s1_address                                (mm_interconnect_0_modo_s1_address),                           //                                  modo_s1.address
		.modo_s1_readdata                               (mm_interconnect_0_modo_s1_readdata),                          //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                         .debugaccess
		.onchip_memory2_0_s1_address                    (mm_interconnect_0_onchip_memory2_0_s1_address),               //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                         .clken
		.push_buttons_s1_address                        (mm_interconnect_0_push_buttons_s1_address),                   //                          push_buttons_s1.address
		.push_buttons_s1_readdata                       (mm_interconnect_0_push_buttons_s1_readdata),                  //                                         .readdata
		.segundos_d_s1_address                          (mm_interconnect_0_segundos_d_s1_address),                     //                            segundos_d_s1.address
		.segundos_d_s1_write                            (mm_interconnect_0_segundos_d_s1_write),                       //                                         .write
		.segundos_d_s1_readdata                         (mm_interconnect_0_segundos_d_s1_readdata),                    //                                         .readdata
		.segundos_d_s1_writedata                        (mm_interconnect_0_segundos_d_s1_writedata),                   //                                         .writedata
		.segundos_d_s1_chipselect                       (mm_interconnect_0_segundos_d_s1_chipselect),                  //                                         .chipselect
		.segundos_u_s1_address                          (mm_interconnect_0_segundos_u_s1_address),                     //                            segundos_u_s1.address
		.segundos_u_s1_write                            (mm_interconnect_0_segundos_u_s1_write),                       //                                         .write
		.segundos_u_s1_readdata                         (mm_interconnect_0_segundos_u_s1_readdata),                    //                                         .readdata
		.segundos_u_s1_writedata                        (mm_interconnect_0_segundos_u_s1_writedata),                   //                                         .writedata
		.segundos_u_s1_chipselect                       (mm_interconnect_0_segundos_u_s1_chipselect),                  //                                         .chipselect
		.timer_0_s1_address                             (mm_interconnect_0_timer_0_s1_address),                        //                               timer_0_s1.address
		.timer_0_s1_write                               (mm_interconnect_0_timer_0_s1_write),                          //                                         .write
		.timer_0_s1_readdata                            (mm_interconnect_0_timer_0_s1_readdata),                       //                                         .readdata
		.timer_0_s1_writedata                           (mm_interconnect_0_timer_0_s1_writedata),                      //                                         .writedata
		.timer_0_s1_chipselect                          (mm_interconnect_0_timer_0_s1_chipselect)                      //                                         .chipselect
	);

	onchipAlarm_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.sender_irq    (nios2_gen2_0_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
